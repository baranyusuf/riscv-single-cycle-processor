module Decoder_5to32 (
    input  [4:0]  IN,
    output reg [31:0] OUT
);
  always @(*) begin
    case (IN)
      5'd0:  OUT = 32'h0000_0001;
      5'd1:  OUT = 32'h0000_0002;
      5'd2:  OUT = 32'h0000_0004;
      5'd3:  OUT = 32'h0000_0008;
      5'd4:  OUT = 32'h0000_0010;
      5'd5:  OUT = 32'h0000_0020;
      5'd6:  OUT = 32'h0000_0040;
      5'd7:  OUT = 32'h0000_0080;
      5'd8:  OUT = 32'h0000_0100;
      5'd9:  OUT = 32'h0000_0200;
      5'd10: OUT = 32'h0000_0400;
      5'd11: OUT = 32'h0000_0800;
      5'd12: OUT = 32'h0000_1000;
      5'd13: OUT = 32'h0000_2000;
      5'd14: OUT = 32'h0000_4000;
      5'd15: OUT = 32'h0000_8000;
      5'd16: OUT = 32'h0001_0000;
      5'd17: OUT = 32'h0002_0000;
      5'd18: OUT = 32'h0004_0000;
      5'd19: OUT = 32'h0008_0000;
      5'd20: OUT = 32'h0010_0000;
      5'd21: OUT = 32'h0020_0000;
      5'd22: OUT = 32'h0040_0000;
      5'd23: OUT = 32'h0080_0000;
      5'd24: OUT = 32'h0100_0000;
      5'd25: OUT = 32'h0200_0000;
      5'd26: OUT = 32'h0400_0000;
      5'd27: OUT = 32'h0800_0000;
      5'd28: OUT = 32'h1000_0000;
      5'd29: OUT = 32'h2000_0000;
      5'd30: OUT = 32'h4000_0000;
      5'd31: OUT = 32'h8000_0000;
      default: OUT = 32'h0000_0000;
    endcase
  end
endmodule